VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO YMG8K16F18L5BR1_Y10_PA_TOP
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN YMG8K16F18L5BR1_Y10_PA_TOP 0 0 ;
  SIZE 685 BY 1230 ;
  SYMMETRY X Y R90 ;
  PIN ADR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 341.87 0.38 342.25 ;
    END
  END ADR[0]
  PIN ADR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 385.91 0.38 386.29 ;
    END
  END ADR[10]
  PIN ADR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 380.42 0.38 380.8 ;
    END
  END ADR[11]
  PIN ADR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 381.1 0.38 381.48 ;
    END
  END ADR[12]
  PIN ADR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 342.9 0.38 343.28 ;
    END
  END ADR[1]
  PIN ADR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 368.61 0.38 368.99 ;
    END
  END ADR[2]
  PIN ADR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 367.71 0.38 368.09 ;
    END
  END ADR[3]
  PIN ADR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 365.63 0.38 366.01 ;
    END
  END ADR[4]
  PIN ADR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 395.7 0.38 396.08 ;
    END
  END ADR[5]
  PIN ADR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 390.48 0.38 390.86 ;
    END
  END ADR[6]
  PIN ADR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 385.23 0.38 385.61 ;
    END
  END ADR[7]
  PIN ADR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 396.38 0.38 396.76 ;
    END
  END ADR[8]
  PIN ADR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 391.16 0.38 391.54 ;
    END
  END ADR[9]
  PIN BUSY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 282.79 0.28 283.07 ;
    END
  END BUSY
  PIN CLEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 259.95 0.38 260.33 ;
    END
  END CLEN
  PIN CLKIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 237.81 0.38 238.19 ;
    END
  END CLKIN
  PIN CS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 305.72 0.38 306.1 ;
    END
  END CS
  PIN DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 325.52 0.38 325.9 ;
    END
  END DIN[0]
  PIN DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 320.12 0.38 320.5 ;
    END
  END DIN[10]
  PIN DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 319.22 0.38 319.6 ;
    END
  END DIN[11]
  PIN DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 213.69 0.38 214.07 ;
    END
  END DIN[12]
  PIN DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 211.89 0.38 212.27 ;
    END
  END DIN[13]
  PIN DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 192.95 0.38 193.33 ;
    END
  END DIN[14]
  PIN DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 194.75 0.38 195.13 ;
    END
  END DIN[15]
  PIN DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 324.62 0.38 325 ;
    END
  END DIN[1]
  PIN DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 321.92 0.38 322.3 ;
    END
  END DIN[2]
  PIN DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 321.02 0.38 321.4 ;
    END
  END DIN[3]
  PIN DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 209.12 0.38 209.5 ;
    END
  END DIN[4]
  PIN DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 214.59 0.38 214.97 ;
    END
  END DIN[5]
  PIN DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 196.55 0.38 196.93 ;
    END
  END DIN[6]
  PIN DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 236.01 0.38 236.39 ;
    END
  END DIN[7]
  PIN DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 323.72 0.38 324.1 ;
    END
  END DIN[8]
  PIN DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 322.82 0.38 323.2 ;
    END
  END DIN[9]
  PIN DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 318.32 0.38 318.7 ;
    END
  END DOUT[0]
  PIN DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 312.92 0.38 313.3 ;
    END
  END DOUT[10]
  PIN DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 312.02 0.38 312.4 ;
    END
  END DOUT[11]
  PIN DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 212.79 0.38 213.17 ;
    END
  END DOUT[12]
  PIN DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 210.99 0.38 211.37 ;
    END
  END DOUT[13]
  PIN DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 193.85 0.38 194.23 ;
    END
  END DOUT[14]
  PIN DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 195.65 0.38 196.03 ;
    END
  END DOUT[15]
  PIN DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 317.42 0.38 317.8 ;
    END
  END DOUT[1]
  PIN DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 314.72 0.38 315.1 ;
    END
  END DOUT[2]
  PIN DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 313.82 0.38 314.2 ;
    END
  END DOUT[3]
  PIN DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 216.95 0.38 217.33 ;
    END
  END DOUT[4]
  PIN DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 308.195 0.38 308.575 ;
    END
  END DOUT[5]
  PIN DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 217.85 0.38 218.23 ;
    END
  END DOUT[6]
  PIN DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 242.22 0.38 242.6 ;
    END
  END DOUT[7]
  PIN DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 316.52 0.38 316.9 ;
    END
  END DOUT[8]
  PIN DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 315.62 0.38 316 ;
    END
  END DOUT[9]
  PIN EEPROM
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 454.15 0.38 454.53 ;
    END
  END EEPROM
  PIN IFREN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 507.97 0.38 508.35 ;
    END
  END IFREN
  PIN ISAVB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 250.65 0.38 251.03 ;
    END
  END ISAVB
  PIN MRGN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 232.41 0.38 232.79 ;
    END
  END MRGN
  PIN READ
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 259.05 0.38 259.43 ;
    END
  END READ
  PIN SRL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 230.61 0.38 230.99 ;
    END
  END SRL
  PIN STATICEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 278.53 0.44 278.97 ;
    END
  END STATICEN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER METAL2 ;
        RECT 39.105 0 49.105 10 ;
    END
    PORT
      LAYER METAL2 ;
        RECT 55.105 0 65.105 10 ;
    END
    PORT
      LAYER METAL2 ;
        RECT 659 0 669 10 ;
    END
    PORT
      LAYER METAL2 ;
        RECT 675 0 685 10 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER METAL2 ;
        RECT 0 0 10 10 ;
    END
    PORT
      LAYER METAL2 ;
        RECT 16 0 26 10 ;
    END
    PORT
      LAYER METAL2 ;
        RECT 627 0 637 10 ;
    END
    PORT
      LAYER METAL2 ;
        RECT 643 0 653 10 ;
    END
  END VSS
  PIN WR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 0 236.91 0.38 237.29 ;
    END
  END WR
  OBS
    LAYER METAL3 ;
      RECT 0 0 685 1230 ;
    LAYER METAL2 ;
      RECT 1 1 684 1229 ;
      RECT 0 507.97 684 508.35 ;
      RECT 0 454.15 684 454.53 ;
      RECT 0 396.38 684 396.76 ;
      RECT 0 395.7 684 396.08 ;
      RECT 0 391.16 684 391.54 ;
      RECT 0 390.48 684 390.86 ;
      RECT 0 385.91 684 386.29 ;
      RECT 0 385.23 684 385.61 ;
      RECT 0 381.1 684 381.48 ;
      RECT 0 380.42 684 380.8 ;
      RECT 0 368.61 684 368.99 ;
      RECT 0 367.71 684 368.09 ;
      RECT 0 365.63 684 366.01 ;
      RECT 0 342.9 684 343.28 ;
      RECT 0 341.87 684 342.25 ;
      RECT 0 325.52 684 325.9 ;
      RECT 0 324.62 684 325 ;
      RECT 0 323.72 684 324.1 ;
      RECT 0 322.82 684 323.2 ;
      RECT 0 321.92 684 322.3 ;
      RECT 0 321.02 684 321.4 ;
      RECT 0 320.12 684 320.5 ;
      RECT 0 319.22 684 319.6 ;
      RECT 0 318.32 684 318.7 ;
      RECT 0 317.42 684 317.8 ;
      RECT 0 316.52 684 316.9 ;
      RECT 0 315.62 684 316 ;
      RECT 0 314.72 684 315.1 ;
      RECT 0 313.82 684 314.2 ;
      RECT 0 312.92 684 313.3 ;
      RECT 0 312.02 684 312.4 ;
      RECT 0 308.195 684 308.575 ;
      RECT 0 305.72 684 306.1 ;
      RECT 0 282.79 684 283.07 ;
      RECT 0 278.53 684 278.97 ;
      RECT 0 259.95 684 260.33 ;
      RECT 0 259.05 684 259.43 ;
      RECT 0 250.65 684 251.03 ;
      RECT 0 242.22 684 242.6 ;
      RECT 0 237.81 684 238.19 ;
      RECT 0 236.91 684 237.29 ;
      RECT 0 236.01 684 236.39 ;
      RECT 0 232.41 684 232.79 ;
      RECT 0 230.61 684 230.99 ;
      RECT 0 217.85 684 218.23 ;
      RECT 0 216.95 684 217.33 ;
      RECT 0 214.59 684 214.97 ;
      RECT 0 213.69 684 214.07 ;
      RECT 0 212.79 684 213.17 ;
      RECT 0 211.89 684 212.27 ;
      RECT 0 210.99 684 211.37 ;
      RECT 0 209.12 684 209.5 ;
      RECT 0 196.55 684 196.93 ;
      RECT 0 195.65 684 196.03 ;
      RECT 0 194.75 684 195.13 ;
      RECT 0 193.85 684 194.23 ;
      RECT 0 192.95 684 193.33 ;
      RECT 675 0 685 10 ;
      RECT 659 0 669 1229 ;
      RECT 643 0 653 1229 ;
      RECT 627 0 637 1229 ;
      RECT 55.105 0 65.105 1229 ;
      RECT 39.105 0 49.105 1229 ;
      RECT 16 0 26 1229 ;
      RECT 0 0 10 10 ;
    LAYER METAL1 ;
      RECT 0 0 685 1230 ;
  END
END YMG8K16F18L5BR1_Y10_PA_TOP

END LIBRARY
